// DESCRIPTION: PlanV Async Fifo SV UVM Testbench
//
// Property of PlanV GmbH, 2024. All rights reserved.
// Licensed under the Solderpad Hardware License, Version 2.0. See the LICENSE file in the project root for more information.
// Contact: yilou.wang@planv.tech

package sv_fifo_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "sv_fifo_sequence_item.svh"
    `include "sv_fifo_sequence.svh"

    `include "sv_fifo_monitor.svh"
    `include "sv_fifo_driver.svh"
    `include "sv_fifo_scoreboard.svh"
    `include "sv_fifo_sequencer.svh"
    `include "sv_fifo_virtual_sequencer.svh"
    `include "sv_fifo_agent.svh"
    `include "sv_fifo_env.svh"

    `include "sv_case_sequence.svh"

    `include "sv_base_test.svh"
    `include "sv_case_test.svh"

endpackage